BZh91AY&SY�uh �߀Rxg����������`�Qsi�u��:Ԁ@ a�i�yM�A�SA�����42h4dɣ��i�0LM4����Hd�jPh  @   ��SA(�jmM�I�i�  ��2dшbi���4�&&�h �	F� F�h�a��)����z���#��4�m�%x|�
4�"�%h�����f� W<W)\}����N��v�̚����<����d�\����)e�j�neH����4x�)QB3q�Ŷ3)KA����<hI�C.X�i�2`Ta2���Ά|B;|��]��y#��S�������,���*s�Н+�/��)Qk��jE�Fư�� 0h-aBIx�A3~m{�4׎�(?Wܦ㿸݄���x�a�tm�mgp�!Cy�����MC�,���jf���Ir܂��!U��`$��?��Ia�]��gE����s  ,��n����A��Dj@4�1��~�;�Z��F�*v��y��ݧS
�D�nِ�G}�4�
���F�1F-��p�M��[�X0޸�=��s�@ųY��쇺��͐/dj��V[^F�����VE6aDZ	@ZT	�4R��V�
KLk ��z��y�J��i� ���P�+��x���:�U4��I�ޓ�v��{���s���m����C!�3��?�������ʡ�sQ ��I�vO�L�w�|ɒ�ݛ]�F�ZG2�Xw�x�*j��T�\w�QAce8���c[lZ��a2T鍕��2¬���e!�,;پ�}���%�Տ���I��������Sw��d����JOߏ�+���M��wf�m�`��P������^��g�oM�!������g:2�x|�`<��33bA����l�yA�̕��K�%���L[țM�BJB���仲׳���ᐊQ}�.��G�����a�%�D�A�}]uy�b�@�P�D���#Q7�����V�ajĎ�.�����G}���1�.��m6n��WlhN�w�2�.q+4*'&x/��"��%�#f=�E��K��,�A��-QGNj�e�=|�ҜԲB���c����
�@� Ɩ0Y�����I�W�!�O��Be�T�H��hbQb�� qq�{8ffz�H.�	 �K��U)z������:a�i��{w,K��Yy��i��S���Z�<̐1@"g$��[�N���z�#j4$"�p�B�1�p��]t�P�G+!y���'�B���Z�:�������{A�I���
�Xr�Ϥ��6)���5�3��Ĥr'#L!��op�V ��Ԧ��[� �Z��>����p�]�P�P��^!}ئ{��q�6ʥ���.����?\LW�ɤƵ��8�H\��a&�i`4�#g/L�B�`bc����^4E�Ӳq�2�<�X1q��0�!��r�E]��v,d]C(�=f�^	��I�!30C�֏7��nF냱 �`��#��A�P=���B��K�cv��ˀz^m���6��xHF��N������=�	��;����}�ƦI��yI$�iA�z���CL��Ős�5�9�$������'C�f`H8���}�CBڍ{���J��@�u9H�*$2�Dl�K��I>&Ń�ɘ^!x�fmr��o�Xj"�B�#P)W^5�BR�kQ��t��"5k��ъA#@������Ե'R5��ECN���m��х�K5R���j6j �`�bRaiRŏ`M��=�Ľ�Y��B��#W�L���-9���H��X��Bh\ˊ�ĳ�"��'2	߅ΰ��+�;	]P���޽�CF���
�&
�0It�	�ܑN$p�Z 